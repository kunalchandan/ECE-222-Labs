-- QD1.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity QD1 is
	port (
		button_pio_export           : in    std_logic_vector(3 downto 0)  := (others => '0'); --           button_pio.export
		clk_clk                     : in    std_logic                     := '0';             --                  clk.clk
		clk_sdram_clk               : out   std_logic;                                        --            clk_sdram.clk
		led_pio_export              : out   std_logic_vector(7 downto 0);                     --              led_pio.export
		reset_reset_n               : in    std_logic                     := '0';             --                reset.reset_n
		sdram_wire_addr             : out   std_logic_vector(11 downto 0);                    --           sdram_wire.addr
		sdram_wire_ba               : out   std_logic_vector(1 downto 0);                     --                     .ba
		sdram_wire_cas_n            : out   std_logic;                                        --                     .cas_n
		sdram_wire_cke              : out   std_logic;                                        --                     .cke
		sdram_wire_cs_n             : out   std_logic;                                        --                     .cs_n
		sdram_wire_dq               : inout std_logic_vector(15 downto 0) := (others => '0'); --                     .dq
		sdram_wire_dqm              : out   std_logic_vector(1 downto 0);                     --                     .dqm
		sdram_wire_ras_n            : out   std_logic;                                        --                     .ras_n
		sdram_wire_we_n             : out   std_logic;                                        --                     .we_n
		switch_pio_export           : in    std_logic_vector(7 downto 0)  := (others => '0'); --           switch_pio.export
		the_altpll_areset_export    : in    std_logic                     := '0';             --    the_altpll_areset.export
		the_altpll_locked_export    : out   std_logic;                                        --    the_altpll_locked.export
		the_altpll_phasedone_export : out   std_logic                                         -- the_altpll_phasedone.export
	);
end entity QD1;

architecture rtl of QD1 is
	component QD1_button_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component QD1_button_pio;

	component QD1_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component QD1_led_pio;

	component QD1_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component QD1_sdram;

	component QD1_switch_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component QD1_switch_pio;

	component QD1_the_altpll is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			c1        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component QD1_the_altpll;

	component QD1_the_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component QD1_the_jtag_uart;

	component QD1_the_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component QD1_the_master;

	component memory_mapped_reset is
		generic (
			ADDR_WIDTH    : integer := 2;
			REGISTER_SIZE : integer := 32
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			avm_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avm_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avm_readdatavalid : out std_logic;                                        -- readdatavalid
			avm_read          : in  std_logic                     := 'X';             -- read
			avm_write         : in  std_logic                     := 'X';             -- write
			avm_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reset_out         : out std_logic                                         -- reset
		);
	end component memory_mapped_reset;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(30 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component QD1_the_onchip_memory2 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component QD1_the_onchip_memory2;

	component orca_timer is
		generic (
			TIMER_WIDTH : integer := 64
		);
		port (
			clk             : in  std_logic                     := 'X';             -- clk
			reset           : in  std_logic                     := 'X';             -- reset
			timer_value     : out std_logic_vector(63 downto 0);                    -- value
			timer_interrupt : out std_logic;                                        -- interrupt
			slave_AWLOCK    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- slave_awlock
			slave_ARCACHE   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_arcache
			slave_ARID      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_arid
			slave_ARLEN     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_arlen
			slave_ARLOCK    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- slave_arlock
			slave_ARSIZE    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- slave_arsize
			slave_ARBURST   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- slave_awburst
			slave_AWBURST   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- slave_awburst
			slave_AWCACHE   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_awcache
			slave_AWID      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_awid
			slave_AWLEN     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_awlen
			slave_AWSIZE    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- slave_awsize
			slave_BID       : out std_logic_vector(3 downto 0);                     -- slave_bid
			slave_RID       : out std_logic_vector(3 downto 0);                     -- slave_rid
			slave_RLAST     : out std_logic;                                        -- slave_rlast
			slave_WID       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- slave_wid
			slave_WLAST     : in  std_logic                     := 'X';             -- slave_wlast
			slave_ARADDR    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- araddr
			slave_ARPROT    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			slave_ARVALID   : in  std_logic                     := 'X';             -- arvalid
			slave_ARREADY   : out std_logic;                                        -- arready
			slave_RDATA     : out std_logic_vector(31 downto 0);                    -- rdata
			slave_RVALID    : out std_logic;                                        -- rvalid
			slave_RREADY    : in  std_logic                     := 'X';             -- rready
			slave_AWADDR    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awaddr
			slave_AWPROT    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			slave_AWVALID   : in  std_logic                     := 'X';             -- awvalid
			slave_AWREADY   : out std_logic;                                        -- awready
			slave_WDATA     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			slave_WSTRB     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			slave_WVALID    : in  std_logic                     := 'X';             -- wvalid
			slave_WREADY    : out std_logic;                                        -- wready
			slave_BVALID    : out std_logic;                                        -- bvalid
			slave_BREADY    : in  std_logic                     := 'X';             -- bready
			slave_BRESP     : out std_logic_vector(1 downto 0);                     -- bresp
			slave_RRESP     : out std_logic_vector(1 downto 0)                      -- rresp
		);
	end component orca_timer;

	component ORCA is
		generic (
			REGISTER_SIZE                : integer                       := 32;
			RESET_VECTOR                 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			ENABLE_EXCEPTIONS            : natural                       := 1;
			INTERRUPT_VECTOR             : std_logic_vector(31 downto 0) := "00000000000000000000001000000000";
			ENABLE_EXT_INTERRUPTS        : natural                       := 1;
			NUM_EXT_INTERRUPTS           : positive                      := 1;
			MAX_IFETCHES_IN_FLIGHT       : natural                       := 1;
			BTB_ENTRIES                  : natural                       := 16;
			MULTIPLY_ENABLE              : natural                       := 1;
			SHIFTER_MAX_CYCLES           : natural                       := 32;
			DIVIDE_ENABLE                : natural                       := 1;
			PIPELINE_STAGES              : natural                       := 4;
			VCP_ENABLE                   : natural                       := 0;
			POWER_OPTIMIZED              : natural                       := 0;
			FAMILY                       : string                        := "INTEL";
			INSTRUCTION_REQUEST_REGISTER : natural                       := 1;
			INSTRUCTION_RETURN_REGISTER  : natural                       := 0;
			DATA_REQUEST_REGISTER        : natural                       := 1;
			DATA_RETURN_REGISTER         : natural                       := 0;
			LOG2_BURSTLENGTH             : positive                      := 4;
			AXI_ID_WIDTH                 : positive                      := 2;
			AVALON_AUX                   : natural                       := 1;
			LMB_AUX                      : natural                       := 0;
			WISHBONE_AUX                 : natural                       := 0;
			ICACHE_SIZE                  : natural                       := 0;
			ICACHE_LINE_SIZE             : natural                       := 32;
			ICACHE_EXTERNAL_WIDTH        : integer                       := 32;
			IC_REQUEST_REGISTER          : natural                       := 1;
			IC_RETURN_REGISTER           : natural                       := 0;
			DCACHE_SIZE                  : natural                       := 0;
			DCACHE_WRITEBACK             : natural                       := 1;
			DCACHE_LINE_SIZE             : natural                       := 32;
			DCACHE_EXTERNAL_WIDTH        : integer                       := 32;
			DC_REQUEST_REGISTER          : natural                       := 1;
			DC_RETURN_REGISTER           : natural                       := 0;
			UC_MEMORY_REGIONS            : natural                       := 0;
			UMR0_ADDR_BASE               : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			UMR0_ADDR_LAST               : std_logic_vector(31 downto 0) := "11111111111111111111111111111111";
			IUC_REQUEST_REGISTER         : natural                       := 0;
			IUC_RETURN_REGISTER          : natural                       := 0;
			DUC_REQUEST_REGISTER         : natural                       := 0;
			DUC_RETURN_REGISTER          : natural                       := 0;
			AUX_MEMORY_REGIONS           : natural                       := 1;
			AMR0_ADDR_BASE               : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			AMR0_ADDR_LAST               : std_logic_vector(31 downto 0) := "11111111111111111111111111111111";
			IAUX_REQUEST_REGISTER        : natural                       := 2;
			IAUX_RETURN_REGISTER         : natural                       := 0;
			DAUX_REQUEST_REGISTER        : natural                       := 2;
			DAUX_RETURN_REGISTER         : natural                       := 0
		);
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			reset                         : in  std_logic                     := 'X';             -- reset
			avm_data_address              : out std_logic_vector(31 downto 0);                    -- address
			avm_data_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_data_read                 : out std_logic;                                        -- read
			avm_data_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_data_write                : out std_logic;                                        -- write
			avm_data_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			avm_data_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			avm_data_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			avm_instruction_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_instruction_read          : out std_logic;                                        -- read
			avm_instruction_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_instruction_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_instruction_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			timer_value                   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- value
			timer_interrupt               : in  std_logic                     := 'X';             -- interrupt
			global_interrupts             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			DUC_ARADDR                    : out std_logic_vector(31 downto 0);                    -- araddr
			DUC_ARBURST                   : out std_logic_vector(1 downto 0);                     -- arburst
			DUC_ARCACHE                   : out std_logic_vector(3 downto 0);                     -- arcache
			DUC_ARID                      : out std_logic_vector(1 downto 0);                     -- arid
			DUC_ARLEN                     : out std_logic_vector(3 downto 0);                     -- arlen
			DUC_ARLOCK                    : out std_logic_vector(1 downto 0);                     -- arlock
			DUC_ARPROT                    : out std_logic_vector(2 downto 0);                     -- arprot
			DUC_ARREADY                   : in  std_logic                     := 'X';             -- arready
			DUC_ARSIZE                    : out std_logic_vector(2 downto 0);                     -- arsize
			DUC_ARVALID                   : out std_logic;                                        -- arvalid
			DUC_AWADDR                    : out std_logic_vector(31 downto 0);                    -- awaddr
			DUC_AWBURST                   : out std_logic_vector(1 downto 0);                     -- awburst
			DUC_AWCACHE                   : out std_logic_vector(3 downto 0);                     -- awcache
			DUC_AWID                      : out std_logic_vector(1 downto 0);                     -- awid
			DUC_AWLEN                     : out std_logic_vector(3 downto 0);                     -- awlen
			DUC_AWLOCK                    : out std_logic_vector(1 downto 0);                     -- awlock
			DUC_AWPROT                    : out std_logic_vector(2 downto 0);                     -- awprot
			DUC_AWREADY                   : in  std_logic                     := 'X';             -- awready
			DUC_AWSIZE                    : out std_logic_vector(2 downto 0);                     -- awsize
			DUC_AWVALID                   : out std_logic;                                        -- awvalid
			DUC_BID                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bid
			DUC_BREADY                    : out std_logic;                                        -- bready
			DUC_BRESP                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			DUC_BVALID                    : in  std_logic                     := 'X';             -- bvalid
			DUC_RDATA                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			DUC_RID                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rid
			DUC_RLAST                     : in  std_logic                     := 'X';             -- rlast
			DUC_RREADY                    : out std_logic;                                        -- rready
			DUC_RRESP                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			DUC_RVALID                    : in  std_logic                     := 'X';             -- rvalid
			DUC_WDATA                     : out std_logic_vector(31 downto 0);                    -- wdata
			DUC_WID                       : out std_logic_vector(1 downto 0);                     -- wid
			DUC_WLAST                     : out std_logic;                                        -- wlast
			DUC_WREADY                    : in  std_logic                     := 'X';             -- wready
			DUC_WSTRB                     : out std_logic_vector(3 downto 0);                     -- wstrb
			DUC_WVALID                    : out std_logic;                                        -- wvalid
			IUC_ARADDR                    : out std_logic_vector(31 downto 0);                    -- araddr
			IUC_ARBURST                   : out std_logic_vector(1 downto 0);                     -- arburst
			IUC_ARCACHE                   : out std_logic_vector(3 downto 0);                     -- arcache
			IUC_ARID                      : out std_logic_vector(1 downto 0);                     -- arid
			IUC_ARLEN                     : out std_logic_vector(3 downto 0);                     -- arlen
			IUC_ARLOCK                    : out std_logic_vector(1 downto 0);                     -- arlock
			IUC_ARPROT                    : out std_logic_vector(2 downto 0);                     -- arprot
			IUC_ARREADY                   : in  std_logic                     := 'X';             -- arready
			IUC_ARSIZE                    : out std_logic_vector(2 downto 0);                     -- arsize
			IUC_ARVALID                   : out std_logic;                                        -- arvalid
			IUC_AWADDR                    : out std_logic_vector(31 downto 0);                    -- awaddr
			IUC_AWBURST                   : out std_logic_vector(1 downto 0);                     -- awburst
			IUC_AWCACHE                   : out std_logic_vector(3 downto 0);                     -- awcache
			IUC_AWID                      : out std_logic_vector(1 downto 0);                     -- awid
			IUC_AWLEN                     : out std_logic_vector(3 downto 0);                     -- awlen
			IUC_AWLOCK                    : out std_logic_vector(1 downto 0);                     -- awlock
			IUC_AWPROT                    : out std_logic_vector(2 downto 0);                     -- awprot
			IUC_AWREADY                   : in  std_logic                     := 'X';             -- awready
			IUC_AWSIZE                    : out std_logic_vector(2 downto 0);                     -- awsize
			IUC_AWVALID                   : out std_logic;                                        -- awvalid
			IUC_BID                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bid
			IUC_BREADY                    : out std_logic;                                        -- bready
			IUC_BRESP                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			IUC_BVALID                    : in  std_logic                     := 'X';             -- bvalid
			IUC_RDATA                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			IUC_RID                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rid
			IUC_RLAST                     : in  std_logic                     := 'X';             -- rlast
			IUC_RREADY                    : out std_logic;                                        -- rready
			IUC_RRESP                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			IUC_RVALID                    : in  std_logic                     := 'X';             -- rvalid
			IUC_WDATA                     : out std_logic_vector(31 downto 0);                    -- wdata
			IUC_WID                       : out std_logic_vector(1 downto 0);                     -- wid
			IUC_WLAST                     : out std_logic;                                        -- wlast
			IUC_WREADY                    : in  std_logic                     := 'X';             -- wready
			IUC_WSTRB                     : out std_logic_vector(3 downto 0);                     -- wstrb
			IUC_WVALID                    : out std_logic;                                        -- wvalid
			IC_ARADDR                     : out std_logic_vector(31 downto 0);                    -- araddr
			IC_ARBURST                    : out std_logic_vector(1 downto 0);                     -- arburst
			IC_ARCACHE                    : out std_logic_vector(3 downto 0);                     -- arcache
			IC_ARID                       : out std_logic_vector(1 downto 0);                     -- arid
			IC_ARLEN                      : out std_logic_vector(3 downto 0);                     -- arlen
			IC_ARLOCK                     : out std_logic_vector(1 downto 0);                     -- arlock
			IC_ARPROT                     : out std_logic_vector(2 downto 0);                     -- arprot
			IC_ARREADY                    : in  std_logic                     := 'X';             -- arready
			IC_ARSIZE                     : out std_logic_vector(2 downto 0);                     -- arsize
			IC_ARVALID                    : out std_logic;                                        -- arvalid
			IC_AWADDR                     : out std_logic_vector(31 downto 0);                    -- awaddr
			IC_AWBURST                    : out std_logic_vector(1 downto 0);                     -- awburst
			IC_AWCACHE                    : out std_logic_vector(3 downto 0);                     -- awcache
			IC_AWID                       : out std_logic_vector(1 downto 0);                     -- awid
			IC_AWLEN                      : out std_logic_vector(3 downto 0);                     -- awlen
			IC_AWLOCK                     : out std_logic_vector(1 downto 0);                     -- awlock
			IC_AWPROT                     : out std_logic_vector(2 downto 0);                     -- awprot
			IC_AWREADY                    : in  std_logic                     := 'X';             -- awready
			IC_AWSIZE                     : out std_logic_vector(2 downto 0);                     -- awsize
			IC_AWVALID                    : out std_logic;                                        -- awvalid
			IC_BID                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bid
			IC_BREADY                     : out std_logic;                                        -- bready
			IC_BRESP                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			IC_BVALID                     : in  std_logic                     := 'X';             -- bvalid
			IC_RDATA                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			IC_RID                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rid
			IC_RLAST                      : in  std_logic                     := 'X';             -- rlast
			IC_RREADY                     : out std_logic;                                        -- rready
			IC_RRESP                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			IC_RVALID                     : in  std_logic                     := 'X';             -- rvalid
			IC_WDATA                      : out std_logic_vector(31 downto 0);                    -- wdata
			IC_WID                        : out std_logic_vector(1 downto 0);                     -- wid
			IC_WLAST                      : out std_logic;                                        -- wlast
			IC_WREADY                     : in  std_logic                     := 'X';             -- wready
			IC_WSTRB                      : out std_logic_vector(3 downto 0);                     -- wstrb
			IC_WVALID                     : out std_logic;                                        -- wvalid
			DC_ARADDR                     : out std_logic_vector(31 downto 0);                    -- araddr
			DC_ARBURST                    : out std_logic_vector(1 downto 0);                     -- arburst
			DC_ARCACHE                    : out std_logic_vector(3 downto 0);                     -- arcache
			DC_ARID                       : out std_logic_vector(1 downto 0);                     -- arid
			DC_ARLEN                      : out std_logic_vector(3 downto 0);                     -- arlen
			DC_ARLOCK                     : out std_logic_vector(1 downto 0);                     -- arlock
			DC_ARPROT                     : out std_logic_vector(2 downto 0);                     -- arprot
			DC_ARREADY                    : in  std_logic                     := 'X';             -- arready
			DC_ARSIZE                     : out std_logic_vector(2 downto 0);                     -- arsize
			DC_ARVALID                    : out std_logic;                                        -- arvalid
			DC_AWADDR                     : out std_logic_vector(31 downto 0);                    -- awaddr
			DC_AWBURST                    : out std_logic_vector(1 downto 0);                     -- awburst
			DC_AWCACHE                    : out std_logic_vector(3 downto 0);                     -- awcache
			DC_AWID                       : out std_logic_vector(1 downto 0);                     -- awid
			DC_AWLEN                      : out std_logic_vector(3 downto 0);                     -- awlen
			DC_AWLOCK                     : out std_logic_vector(1 downto 0);                     -- awlock
			DC_AWPROT                     : out std_logic_vector(2 downto 0);                     -- awprot
			DC_AWREADY                    : in  std_logic                     := 'X';             -- awready
			DC_AWSIZE                     : out std_logic_vector(2 downto 0);                     -- awsize
			DC_AWVALID                    : out std_logic;                                        -- awvalid
			DC_BID                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bid
			DC_BREADY                     : out std_logic;                                        -- bready
			DC_BRESP                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			DC_BVALID                     : in  std_logic                     := 'X';             -- bvalid
			DC_RDATA                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			DC_RID                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rid
			DC_RLAST                      : in  std_logic                     := 'X';             -- rlast
			DC_RREADY                     : out std_logic;                                        -- rready
			DC_RRESP                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			DC_RVALID                     : in  std_logic                     := 'X';             -- rvalid
			DC_WDATA                      : out std_logic_vector(31 downto 0);                    -- wdata
			DC_WID                        : out std_logic_vector(1 downto 0);                     -- wid
			DC_WLAST                      : out std_logic;                                        -- wlast
			DC_WREADY                     : in  std_logic                     := 'X';             -- wready
			DC_WSTRB                      : out std_logic_vector(3 downto 0);                     -- wstrb
			DC_WVALID                     : out std_logic;                                        -- wvalid
			vcp_data0                     : out std_logic_vector(31 downto 0);                    -- data0
			vcp_data1                     : out std_logic_vector(31 downto 0);                    -- data1
			vcp_data2                     : out std_logic_vector(31 downto 0);                    -- data2
			vcp_instruction               : out std_logic_vector(40 downto 0);                    -- instruction
			vcp_valid_instr               : out std_logic;                                        -- valid_instr
			vcp_ready                     : in  std_logic                     := 'X';             -- ready
			vcp_illegal                   : in  std_logic                     := 'X';             -- illegal
			vcp_writeback_data            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writeback_data
			vcp_writeback_en              : in  std_logic                     := 'X';             -- writeback_en
			vcp_alu_data1                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- alu_data1
			vcp_alu_data2                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- alu_data2
			vcp_alu_source_valid          : in  std_logic                     := 'X';             -- alu_source_valid
			vcp_alu_result                : out std_logic_vector(31 downto 0);                    -- alu_result
			vcp_alu_result_valid          : out std_logic;                                        -- alu_result_valid
			data_ADR_O                    : out std_logic_vector(31 downto 0);                    -- ADR_O
			data_DAT_I                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DAT_I
			data_DAT_O                    : out std_logic_vector(31 downto 0);                    -- DAT_O
			data_WE_O                     : out std_logic;                                        -- WE_O
			data_SEL_O                    : out std_logic_vector(3 downto 0);                     -- SEL_O
			data_STB_O                    : out std_logic;                                        -- STB_O
			data_ACK_I                    : in  std_logic                     := 'X';             -- ACK_I
			data_CYC_O                    : out std_logic;                                        -- CYC_O
			data_CTI_O                    : out std_logic_vector(2 downto 0);                     -- CTI_O
			data_STALL_I                  : in  std_logic                     := 'X';             -- STALL_I
			instr_ADR_O                   : out std_logic_vector(31 downto 0);                    -- ADR_O
			instr_DAT_I                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DAT_I
			instr_STB_O                   : out std_logic;                                        -- STB_O
			instr_ACK_I                   : in  std_logic                     := 'X';             -- ACK_I
			instr_CYC_O                   : out std_logic;                                        -- CYC_O
			instr_CTI_O                   : out std_logic_vector(2 downto 0);                     -- CTI_O
			instr_STALL_I                 : in  std_logic                     := 'X';             -- STALL_I
			ILMB_Addr                     : out std_logic_vector(31 downto 0);                    -- Addr
			ILMB_Byte_Enable              : out std_logic_vector(3 downto 0);                     -- Byte_Enable
			ILMB_Data_Write               : out std_logic_vector(31 downto 0);                    -- Data_Write
			ILMB_AS                       : out std_logic;                                        -- AS
			ILMB_Read_Strobe              : out std_logic;                                        -- Read_Strobe
			ILMB_Write_Strobe             : out std_logic;                                        -- Write_Strobe
			ILMB_Data_Read                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- Data_Read
			ILMB_Ready                    : in  std_logic                     := 'X';             -- Ready
			ILMB_Wait                     : in  std_logic                     := 'X';             -- Wait
			ILMB_CE                       : in  std_logic                     := 'X';             -- CE
			ILMB_UE                       : in  std_logic                     := 'X';             -- UE
			DLMB_Addr                     : out std_logic_vector(31 downto 0);                    -- Addr
			DLMB_Byte_Enable              : out std_logic_vector(3 downto 0);                     -- Byte_Enable
			DLMB_Data_Write               : out std_logic_vector(31 downto 0);                    -- Data_Write
			DLMB_AS                       : out std_logic;                                        -- AS
			DLMB_Read_Strobe              : out std_logic;                                        -- Read_Strobe
			DLMB_Write_Strobe             : out std_logic;                                        -- Write_Strobe
			DLMB_Data_Read                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- Data_Read
			DLMB_Ready                    : in  std_logic                     := 'X';             -- Ready
			DLMB_Wait                     : in  std_logic                     := 'X';             -- Wait
			DLMB_CE                       : in  std_logic                     := 'X';             -- CE
			DLMB_UE                       : in  std_logic                     := 'X'              -- UE
		);
	end component ORCA;

	component QD1_mm_interconnect_0 is
		port (
			the_orca_timer_slave_awaddr                                       : out std_logic_vector(3 downto 0);                     -- awaddr
			the_orca_timer_slave_awprot                                       : out std_logic_vector(2 downto 0);                     -- awprot
			the_orca_timer_slave_awvalid                                      : out std_logic;                                        -- awvalid
			the_orca_timer_slave_awready                                      : in  std_logic                     := 'X';             -- awready
			the_orca_timer_slave_wdata                                        : out std_logic_vector(31 downto 0);                    -- wdata
			the_orca_timer_slave_wstrb                                        : out std_logic_vector(3 downto 0);                     -- wstrb
			the_orca_timer_slave_wvalid                                       : out std_logic;                                        -- wvalid
			the_orca_timer_slave_wready                                       : in  std_logic                     := 'X';             -- wready
			the_orca_timer_slave_bresp                                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			the_orca_timer_slave_bvalid                                       : in  std_logic                     := 'X';             -- bvalid
			the_orca_timer_slave_bready                                       : out std_logic;                                        -- bready
			the_orca_timer_slave_araddr                                       : out std_logic_vector(3 downto 0);                     -- araddr
			the_orca_timer_slave_arprot                                       : out std_logic_vector(2 downto 0);                     -- arprot
			the_orca_timer_slave_arvalid                                      : out std_logic;                                        -- arvalid
			the_orca_timer_slave_arready                                      : in  std_logic                     := 'X';             -- arready
			the_orca_timer_slave_rdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			the_orca_timer_slave_rresp                                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			the_orca_timer_slave_rvalid                                       : in  std_logic                     := 'X';             -- rvalid
			the_orca_timer_slave_rready                                       : out std_logic;                                        -- rready
			the_altpll_c0_clk                                                 : in  std_logic                     := 'X';             -- clk
			the_clk_clk_clk                                                   : in  std_logic                     := 'X';             -- clk
			the_altpll_inclk_interface_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			the_jtag_uart_reset_reset_bridge_in_reset_reset                   : in  std_logic                     := 'X';             -- reset
			the_master_clk_reset_reset_bridge_in_reset_reset                  : in  std_logic                     := 'X';             -- reset
			the_mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			the_vectorblox_orca_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			the_master_master_address                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			the_master_master_waitrequest                                     : out std_logic;                                        -- waitrequest
			the_master_master_byteenable                                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			the_master_master_read                                            : in  std_logic                     := 'X';             -- read
			the_master_master_readdata                                        : out std_logic_vector(31 downto 0);                    -- readdata
			the_master_master_readdatavalid                                   : out std_logic;                                        -- readdatavalid
			the_master_master_write                                           : in  std_logic                     := 'X';             -- write
			the_master_master_writedata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			the_mm_clock_crossing_bridge_m0_address                           : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			the_mm_clock_crossing_bridge_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			the_mm_clock_crossing_bridge_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			the_mm_clock_crossing_bridge_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			the_mm_clock_crossing_bridge_m0_read                              : in  std_logic                     := 'X';             -- read
			the_mm_clock_crossing_bridge_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			the_mm_clock_crossing_bridge_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			the_mm_clock_crossing_bridge_m0_write                             : in  std_logic                     := 'X';             -- write
			the_mm_clock_crossing_bridge_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			the_mm_clock_crossing_bridge_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			the_vectorblox_orca_data_address                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			the_vectorblox_orca_data_waitrequest                              : out std_logic;                                        -- waitrequest
			the_vectorblox_orca_data_byteenable                               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			the_vectorblox_orca_data_read                                     : in  std_logic                     := 'X';             -- read
			the_vectorblox_orca_data_readdata                                 : out std_logic_vector(31 downto 0);                    -- readdata
			the_vectorblox_orca_data_readdatavalid                            : out std_logic;                                        -- readdatavalid
			the_vectorblox_orca_data_write                                    : in  std_logic                     := 'X';             -- write
			the_vectorblox_orca_data_writedata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			button_pio_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			button_pio_s1_write                                               : out std_logic;                                        -- write
			button_pio_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_pio_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			button_pio_s1_chipselect                                          : out std_logic;                                        -- chipselect
			led_pio_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                                                  : out std_logic;                                        -- write
			led_pio_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                                             : out std_logic;                                        -- chipselect
			sdram_s1_address                                                  : out std_logic_vector(21 downto 0);                    -- address
			sdram_s1_write                                                    : out std_logic;                                        -- write
			sdram_s1_read                                                     : out std_logic;                                        -- read
			sdram_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                               : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                            : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                              : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                               : out std_logic;                                        -- chipselect
			switch_pio_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			switch_pio_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_altpll_pll_slave_address                                      : out std_logic_vector(1 downto 0);                     -- address
			the_altpll_pll_slave_write                                        : out std_logic;                                        -- write
			the_altpll_pll_slave_read                                         : out std_logic;                                        -- read
			the_altpll_pll_slave_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_altpll_pll_slave_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			the_jtag_uart_avalon_jtag_slave_address                           : out std_logic_vector(0 downto 0);                     -- address
			the_jtag_uart_avalon_jtag_slave_write                             : out std_logic;                                        -- write
			the_jtag_uart_avalon_jtag_slave_read                              : out std_logic;                                        -- read
			the_jtag_uart_avalon_jtag_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_jtag_uart_avalon_jtag_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			the_jtag_uart_avalon_jtag_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			the_jtag_uart_avalon_jtag_slave_chipselect                        : out std_logic;                                        -- chipselect
			the_memory_mapped_reset_avalon_slave_address                      : out std_logic_vector(1 downto 0);                     -- address
			the_memory_mapped_reset_avalon_slave_write                        : out std_logic;                                        -- write
			the_memory_mapped_reset_avalon_slave_read                         : out std_logic;                                        -- read
			the_memory_mapped_reset_avalon_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_memory_mapped_reset_avalon_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			the_memory_mapped_reset_avalon_slave_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			the_mm_clock_crossing_bridge_s0_address                           : out std_logic_vector(30 downto 0);                    -- address
			the_mm_clock_crossing_bridge_s0_write                             : out std_logic;                                        -- write
			the_mm_clock_crossing_bridge_s0_read                              : out std_logic;                                        -- read
			the_mm_clock_crossing_bridge_s0_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_mm_clock_crossing_bridge_s0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			the_mm_clock_crossing_bridge_s0_burstcount                        : out std_logic_vector(0 downto 0);                     -- burstcount
			the_mm_clock_crossing_bridge_s0_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			the_mm_clock_crossing_bridge_s0_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			the_mm_clock_crossing_bridge_s0_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			the_mm_clock_crossing_bridge_s0_debugaccess                       : out std_logic;                                        -- debugaccess
			the_onchip_memory2_s2_address                                     : out std_logic_vector(12 downto 0);                    -- address
			the_onchip_memory2_s2_write                                       : out std_logic;                                        -- write
			the_onchip_memory2_s2_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_onchip_memory2_s2_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			the_onchip_memory2_s2_byteenable                                  : out std_logic_vector(3 downto 0);                     -- byteenable
			the_onchip_memory2_s2_chipselect                                  : out std_logic;                                        -- chipselect
			the_onchip_memory2_s2_clken                                       : out std_logic                                         -- clken
		);
	end component QD1_mm_interconnect_0;

	component QD1_mm_interconnect_1 is
		port (
			the_altpll_c0_clk                                     : in  std_logic                     := 'X';             -- clk
			the_onchip_memory2_reset1_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			the_vectorblox_orca_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			the_vectorblox_orca_instruction_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			the_vectorblox_orca_instruction_waitrequest           : out std_logic;                                        -- waitrequest
			the_vectorblox_orca_instruction_read                  : in  std_logic                     := 'X';             -- read
			the_vectorblox_orca_instruction_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			the_vectorblox_orca_instruction_readdatavalid         : out std_logic;                                        -- readdatavalid
			the_onchip_memory2_s1_address                         : out std_logic_vector(12 downto 0);                    -- address
			the_onchip_memory2_s1_write                           : out std_logic;                                        -- write
			the_onchip_memory2_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			the_onchip_memory2_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			the_onchip_memory2_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			the_onchip_memory2_s1_chipselect                      : out std_logic;                                        -- chipselect
			the_onchip_memory2_s1_clken                           : out std_logic                                         -- clken
		);
	end component QD1_mm_interconnect_1;

	component QD1_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component QD1_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component qd1_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component qd1_rst_controller;

	component qd1_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component qd1_rst_controller_001;

	component qd1_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component qd1_rst_controller_002;

	signal the_altpll_c0_clk                                                    : std_logic;                     -- the_altpll:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, mm_interconnect_0:the_altpll_c0_clk, mm_interconnect_1:the_altpll_c0_clk, rst_controller_001:clk, rst_controller_003:clk, sdram:clk, the_mm_clock_crossing_bridge:s0_clk, the_onchip_memory2:clk, the_onchip_memory2:clk2, the_orca_timer:clk, the_vectorblox_orca:clk]
	signal the_orca_timer_timer_interface_interrupt                             : std_logic;                     -- the_orca_timer:timer_interrupt -> the_vectorblox_orca:timer_interrupt
	signal the_orca_timer_timer_interface_value                                 : std_logic_vector(63 downto 0); -- the_orca_timer:timer_value -> the_vectorblox_orca:timer_value
	signal the_vectorblox_orca_data_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_vectorblox_orca_data_readdata -> the_vectorblox_orca:avm_data_readdata
	signal the_vectorblox_orca_data_waitrequest                                 : std_logic;                     -- mm_interconnect_0:the_vectorblox_orca_data_waitrequest -> the_vectorblox_orca:avm_data_waitrequest
	signal the_vectorblox_orca_data_address                                     : std_logic_vector(31 downto 0); -- the_vectorblox_orca:avm_data_address -> mm_interconnect_0:the_vectorblox_orca_data_address
	signal the_vectorblox_orca_data_byteenable                                  : std_logic_vector(3 downto 0);  -- the_vectorblox_orca:avm_data_byteenable -> mm_interconnect_0:the_vectorblox_orca_data_byteenable
	signal the_vectorblox_orca_data_read                                        : std_logic;                     -- the_vectorblox_orca:avm_data_read -> mm_interconnect_0:the_vectorblox_orca_data_read
	signal the_vectorblox_orca_data_readdatavalid                               : std_logic;                     -- mm_interconnect_0:the_vectorblox_orca_data_readdatavalid -> the_vectorblox_orca:avm_data_readdatavalid
	signal the_vectorblox_orca_data_write                                       : std_logic;                     -- the_vectorblox_orca:avm_data_write -> mm_interconnect_0:the_vectorblox_orca_data_write
	signal the_vectorblox_orca_data_writedata                                   : std_logic_vector(31 downto 0); -- the_vectorblox_orca:avm_data_writedata -> mm_interconnect_0:the_vectorblox_orca_data_writedata
	signal the_master_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_master_master_readdata -> the_master:master_readdata
	signal the_master_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:the_master_master_waitrequest -> the_master:master_waitrequest
	signal the_master_master_address                                            : std_logic_vector(31 downto 0); -- the_master:master_address -> mm_interconnect_0:the_master_master_address
	signal the_master_master_read                                               : std_logic;                     -- the_master:master_read -> mm_interconnect_0:the_master_master_read
	signal the_master_master_byteenable                                         : std_logic_vector(3 downto 0);  -- the_master:master_byteenable -> mm_interconnect_0:the_master_master_byteenable
	signal the_master_master_readdatavalid                                      : std_logic;                     -- mm_interconnect_0:the_master_master_readdatavalid -> the_master:master_readdatavalid
	signal the_master_master_write                                              : std_logic;                     -- the_master:master_write -> mm_interconnect_0:the_master_master_write
	signal the_master_master_writedata                                          : std_logic_vector(31 downto 0); -- the_master:master_writedata -> mm_interconnect_0:the_master_master_writedata
	signal the_mm_clock_crossing_bridge_m0_waitrequest                          : std_logic;                     -- mm_interconnect_0:the_mm_clock_crossing_bridge_m0_waitrequest -> the_mm_clock_crossing_bridge:m0_waitrequest
	signal the_mm_clock_crossing_bridge_m0_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_mm_clock_crossing_bridge_m0_readdata -> the_mm_clock_crossing_bridge:m0_readdata
	signal the_mm_clock_crossing_bridge_m0_debugaccess                          : std_logic;                     -- the_mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_debugaccess
	signal the_mm_clock_crossing_bridge_m0_address                              : std_logic_vector(30 downto 0); -- the_mm_clock_crossing_bridge:m0_address -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_address
	signal the_mm_clock_crossing_bridge_m0_read                                 : std_logic;                     -- the_mm_clock_crossing_bridge:m0_read -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_read
	signal the_mm_clock_crossing_bridge_m0_byteenable                           : std_logic_vector(3 downto 0);  -- the_mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_byteenable
	signal the_mm_clock_crossing_bridge_m0_readdatavalid                        : std_logic;                     -- mm_interconnect_0:the_mm_clock_crossing_bridge_m0_readdatavalid -> the_mm_clock_crossing_bridge:m0_readdatavalid
	signal the_mm_clock_crossing_bridge_m0_writedata                            : std_logic_vector(31 downto 0); -- the_mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_writedata
	signal the_mm_clock_crossing_bridge_m0_write                                : std_logic;                     -- the_mm_clock_crossing_bridge:m0_write -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_write
	signal the_mm_clock_crossing_bridge_m0_burstcount                           : std_logic_vector(0 downto 0);  -- the_mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_0:the_mm_clock_crossing_bridge_m0_burstcount
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_readdata           : std_logic_vector(31 downto 0); -- the_mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:the_mm_clock_crossing_bridge_s0_readdata
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_waitrequest        : std_logic;                     -- the_mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:the_mm_clock_crossing_bridge_s0_waitrequest
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_debugaccess        : std_logic;                     -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_debugaccess -> the_mm_clock_crossing_bridge:s0_debugaccess
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_address            : std_logic_vector(30 downto 0); -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_address -> the_mm_clock_crossing_bridge:s0_address
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_read               : std_logic;                     -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_read -> the_mm_clock_crossing_bridge:s0_read
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_byteenable -> the_mm_clock_crossing_bridge:s0_byteenable
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_readdatavalid      : std_logic;                     -- the_mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:the_mm_clock_crossing_bridge_s0_readdatavalid
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_write              : std_logic;                     -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_write -> the_mm_clock_crossing_bridge:s0_write
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_writedata -> the_mm_clock_crossing_bridge:s0_writedata
	signal mm_interconnect_0_the_mm_clock_crossing_bridge_s0_burstcount         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:the_mm_clock_crossing_bridge_s0_burstcount -> the_mm_clock_crossing_bridge:s0_burstcount
	signal mm_interconnect_0_the_onchip_memory2_s2_chipselect                   : std_logic;                     -- mm_interconnect_0:the_onchip_memory2_s2_chipselect -> the_onchip_memory2:chipselect2
	signal mm_interconnect_0_the_onchip_memory2_s2_readdata                     : std_logic_vector(31 downto 0); -- the_onchip_memory2:readdata2 -> mm_interconnect_0:the_onchip_memory2_s2_readdata
	signal mm_interconnect_0_the_onchip_memory2_s2_address                      : std_logic_vector(12 downto 0); -- mm_interconnect_0:the_onchip_memory2_s2_address -> the_onchip_memory2:address2
	signal mm_interconnect_0_the_onchip_memory2_s2_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:the_onchip_memory2_s2_byteenable -> the_onchip_memory2:byteenable2
	signal mm_interconnect_0_the_onchip_memory2_s2_write                        : std_logic;                     -- mm_interconnect_0:the_onchip_memory2_s2_write -> the_onchip_memory2:write2
	signal mm_interconnect_0_the_onchip_memory2_s2_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_onchip_memory2_s2_writedata -> the_onchip_memory2:writedata2
	signal mm_interconnect_0_the_onchip_memory2_s2_clken                        : std_logic;                     -- mm_interconnect_0:the_onchip_memory2_s2_clken -> the_onchip_memory2:clken2
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_chipselect         : std_logic;                     -- mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_chipselect -> the_jtag_uart:av_chipselect
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_readdata           : std_logic_vector(31 downto 0); -- the_jtag_uart:av_readdata -> mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_waitrequest        : std_logic;                     -- the_jtag_uart:av_waitrequest -> mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_address -> the_jtag_uart:av_address
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read               : std_logic;                     -- mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write              : std_logic;                     -- mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_jtag_uart_avalon_jtag_slave_writedata -> the_jtag_uart:av_writedata
	signal mm_interconnect_0_the_memory_mapped_reset_avalon_slave_readdata      : std_logic_vector(31 downto 0); -- the_memory_mapped_reset:avm_readdata -> mm_interconnect_0:the_memory_mapped_reset_avalon_slave_readdata
	signal mm_interconnect_0_the_memory_mapped_reset_avalon_slave_address       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:the_memory_mapped_reset_avalon_slave_address -> the_memory_mapped_reset:avm_address
	signal mm_interconnect_0_the_memory_mapped_reset_avalon_slave_read          : std_logic;                     -- mm_interconnect_0:the_memory_mapped_reset_avalon_slave_read -> the_memory_mapped_reset:avm_read
	signal mm_interconnect_0_the_memory_mapped_reset_avalon_slave_readdatavalid : std_logic;                     -- the_memory_mapped_reset:avm_readdatavalid -> mm_interconnect_0:the_memory_mapped_reset_avalon_slave_readdatavalid
	signal mm_interconnect_0_the_memory_mapped_reset_avalon_slave_write         : std_logic;                     -- mm_interconnect_0:the_memory_mapped_reset_avalon_slave_write -> the_memory_mapped_reset:avm_write
	signal mm_interconnect_0_the_memory_mapped_reset_avalon_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_memory_mapped_reset_avalon_slave_writedata -> the_memory_mapped_reset:avm_writedata
	signal mm_interconnect_0_the_altpll_pll_slave_readdata                      : std_logic_vector(31 downto 0); -- the_altpll:readdata -> mm_interconnect_0:the_altpll_pll_slave_readdata
	signal mm_interconnect_0_the_altpll_pll_slave_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:the_altpll_pll_slave_address -> the_altpll:address
	signal mm_interconnect_0_the_altpll_pll_slave_read                          : std_logic;                     -- mm_interconnect_0:the_altpll_pll_slave_read -> the_altpll:read
	signal mm_interconnect_0_the_altpll_pll_slave_write                         : std_logic;                     -- mm_interconnect_0:the_altpll_pll_slave_write -> the_altpll:write
	signal mm_interconnect_0_the_altpll_pll_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_altpll_pll_slave_writedata -> the_altpll:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                  : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                               : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                   : std_logic_vector(21 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                      : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                             : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                     : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_led_pio_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                                : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_write                                   : std_logic;                     -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_0_button_pio_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	signal mm_interconnect_0_button_pio_s1_readdata                             : std_logic_vector(31 downto 0); -- button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	signal mm_interconnect_0_button_pio_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_pio_s1_address -> button_pio:address
	signal mm_interconnect_0_button_pio_s1_write                                : std_logic;                     -- mm_interconnect_0:button_pio_s1_write -> mm_interconnect_0_button_pio_s1_write:in
	signal mm_interconnect_0_button_pio_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	signal mm_interconnect_0_switch_pio_s1_readdata                             : std_logic_vector(31 downto 0); -- switch_pio:readdata -> mm_interconnect_0:switch_pio_s1_readdata
	signal mm_interconnect_0_switch_pio_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_pio_s1_address -> switch_pio:address
	signal mm_interconnect_0_the_orca_timer_slave_awaddr                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:the_orca_timer_slave_awaddr -> the_orca_timer:slave_AWADDR
	signal mm_interconnect_0_the_orca_timer_slave_bresp                         : std_logic_vector(1 downto 0);  -- the_orca_timer:slave_BRESP -> mm_interconnect_0:the_orca_timer_slave_bresp
	signal mm_interconnect_0_the_orca_timer_slave_arready                       : std_logic;                     -- the_orca_timer:slave_ARREADY -> mm_interconnect_0:the_orca_timer_slave_arready
	signal mm_interconnect_0_the_orca_timer_slave_rdata                         : std_logic_vector(31 downto 0); -- the_orca_timer:slave_RDATA -> mm_interconnect_0:the_orca_timer_slave_rdata
	signal mm_interconnect_0_the_orca_timer_slave_wstrb                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:the_orca_timer_slave_wstrb -> the_orca_timer:slave_WSTRB
	signal mm_interconnect_0_the_orca_timer_slave_wready                        : std_logic;                     -- the_orca_timer:slave_WREADY -> mm_interconnect_0:the_orca_timer_slave_wready
	signal mm_interconnect_0_the_orca_timer_slave_awready                       : std_logic;                     -- the_orca_timer:slave_AWREADY -> mm_interconnect_0:the_orca_timer_slave_awready
	signal mm_interconnect_0_the_orca_timer_slave_rready                        : std_logic;                     -- mm_interconnect_0:the_orca_timer_slave_rready -> the_orca_timer:slave_RREADY
	signal mm_interconnect_0_the_orca_timer_slave_bready                        : std_logic;                     -- mm_interconnect_0:the_orca_timer_slave_bready -> the_orca_timer:slave_BREADY
	signal mm_interconnect_0_the_orca_timer_slave_wvalid                        : std_logic;                     -- mm_interconnect_0:the_orca_timer_slave_wvalid -> the_orca_timer:slave_WVALID
	signal mm_interconnect_0_the_orca_timer_slave_araddr                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:the_orca_timer_slave_araddr -> the_orca_timer:slave_ARADDR
	signal mm_interconnect_0_the_orca_timer_slave_arprot                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:the_orca_timer_slave_arprot -> the_orca_timer:slave_ARPROT
	signal mm_interconnect_0_the_orca_timer_slave_rresp                         : std_logic_vector(1 downto 0);  -- the_orca_timer:slave_RRESP -> mm_interconnect_0:the_orca_timer_slave_rresp
	signal mm_interconnect_0_the_orca_timer_slave_awprot                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:the_orca_timer_slave_awprot -> the_orca_timer:slave_AWPROT
	signal mm_interconnect_0_the_orca_timer_slave_wdata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:the_orca_timer_slave_wdata -> the_orca_timer:slave_WDATA
	signal mm_interconnect_0_the_orca_timer_slave_arvalid                       : std_logic;                     -- mm_interconnect_0:the_orca_timer_slave_arvalid -> the_orca_timer:slave_ARVALID
	signal mm_interconnect_0_the_orca_timer_slave_bvalid                        : std_logic;                     -- the_orca_timer:slave_BVALID -> mm_interconnect_0:the_orca_timer_slave_bvalid
	signal mm_interconnect_0_the_orca_timer_slave_awvalid                       : std_logic;                     -- mm_interconnect_0:the_orca_timer_slave_awvalid -> the_orca_timer:slave_AWVALID
	signal mm_interconnect_0_the_orca_timer_slave_rvalid                        : std_logic;                     -- the_orca_timer:slave_RVALID -> mm_interconnect_0:the_orca_timer_slave_rvalid
	signal the_vectorblox_orca_instruction_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_1:the_vectorblox_orca_instruction_readdata -> the_vectorblox_orca:avm_instruction_readdata
	signal the_vectorblox_orca_instruction_waitrequest                          : std_logic;                     -- mm_interconnect_1:the_vectorblox_orca_instruction_waitrequest -> the_vectorblox_orca:avm_instruction_waitrequest
	signal the_vectorblox_orca_instruction_address                              : std_logic_vector(31 downto 0); -- the_vectorblox_orca:avm_instruction_address -> mm_interconnect_1:the_vectorblox_orca_instruction_address
	signal the_vectorblox_orca_instruction_read                                 : std_logic;                     -- the_vectorblox_orca:avm_instruction_read -> mm_interconnect_1:the_vectorblox_orca_instruction_read
	signal the_vectorblox_orca_instruction_readdatavalid                        : std_logic;                     -- mm_interconnect_1:the_vectorblox_orca_instruction_readdatavalid -> the_vectorblox_orca:avm_instruction_readdatavalid
	signal mm_interconnect_1_the_onchip_memory2_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:the_onchip_memory2_s1_chipselect -> the_onchip_memory2:chipselect
	signal mm_interconnect_1_the_onchip_memory2_s1_readdata                     : std_logic_vector(31 downto 0); -- the_onchip_memory2:readdata -> mm_interconnect_1:the_onchip_memory2_s1_readdata
	signal mm_interconnect_1_the_onchip_memory2_s1_address                      : std_logic_vector(12 downto 0); -- mm_interconnect_1:the_onchip_memory2_s1_address -> the_onchip_memory2:address
	signal mm_interconnect_1_the_onchip_memory2_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_1:the_onchip_memory2_s1_byteenable -> the_onchip_memory2:byteenable
	signal mm_interconnect_1_the_onchip_memory2_s1_write                        : std_logic;                     -- mm_interconnect_1:the_onchip_memory2_s1_write -> the_onchip_memory2:write
	signal mm_interconnect_1_the_onchip_memory2_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:the_onchip_memory2_s1_writedata -> the_onchip_memory2:writedata
	signal mm_interconnect_1_the_onchip_memory2_s1_clken                        : std_logic;                     -- mm_interconnect_1:the_onchip_memory2_s1_clken -> the_onchip_memory2:clken
	signal the_vectorblox_orca_global_interrupts_irq                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> the_vectorblox_orca:global_interrupts
	signal irq_mapper_receiver0_irq                                             : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                        : std_logic_vector(0 downto 0);  -- the_jtag_uart:av_irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                             : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                                    : std_logic_vector(0 downto 0);  -- button_pio:irq -> irq_synchronizer_001:receiver_irq
	signal rst_controller_reset_out_reset                                       : std_logic;                     -- rst_controller:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_0:the_jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal the_memory_mapped_reset_reset_source_reset                           : std_logic;                     -- the_memory_mapped_reset:reset_out -> [rst_controller:reset_in1, rst_controller_003:reset_in1]
	signal rst_controller_001_reset_out_reset                                   : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:the_mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:the_onchip_memory2_reset1_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset, the_mm_clock_crossing_bridge:s0_reset, the_onchip_memory2:reset, the_onchip_memory2:reset2, the_orca_timer:reset]
	signal rst_controller_001_reset_out_reset_req                               : std_logic;                     -- rst_controller_001:reset_req -> [rst_translator:reset_req_in, the_onchip_memory2:reset_req, the_onchip_memory2:reset_req2]
	signal rst_controller_002_reset_out_reset                                   : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:the_altpll_inclk_interface_reset_reset_bridge_in_reset_reset, mm_interconnect_0:the_master_clk_reset_reset_bridge_in_reset_reset, the_altpll:reset, the_memory_mapped_reset:reset, the_mm_clock_crossing_bridge:m0_reset]
	signal rst_controller_003_reset_out_reset                                   : std_logic;                     -- rst_controller_003:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:the_vectorblox_orca_reset_reset_bridge_in_reset_reset, mm_interconnect_1:the_vectorblox_orca_reset_reset_bridge_in_reset_reset, the_vectorblox_orca:reset]
	signal reset_reset_n_ports_inv                                              : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, the_master:clk_reset_reset]
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read_ports_inv     : std_logic;                     -- mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read:inv -> the_jtag_uart:av_read_n
	signal mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write_ports_inv    : std_logic;                     -- mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write:inv -> the_jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                            : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_0_button_pio_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_button_pio_s1_write:inv -> button_pio:write_n
	signal rst_controller_reset_out_reset_ports_inv                             : std_logic;                     -- rst_controller_reset_out_reset:inv -> [button_pio:reset_n, led_pio:reset_n, switch_pio:reset_n, the_jtag_uart:rst_n]
	signal rst_controller_001_reset_out_reset_ports_inv                         : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> sdram:reset_n

begin

	button_pio : component QD1_button_pio
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_button_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_pio_s1_readdata,        --                    .readdata
			in_port    => button_pio_export,                               -- external_connection.export
			irq        => irq_synchronizer_001_receiver_irq(0)             --                 irq.irq
		);

	led_pio : component QD1_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_export                                -- external_connection.export
		);

	sdram : component QD1_sdram
		port map (
			clk            => the_altpll_c0_clk,                               --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	switch_pio : component QD1_switch_pio
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_switch_pio_s1_readdata, --                    .readdata
			in_port  => switch_pio_export                         -- external_connection.export
		);

	the_altpll : component QD1_the_altpll
		port map (
			clk       => clk_clk,                                          --       inclk_interface.clk
			reset     => rst_controller_002_reset_out_reset,               -- inclk_interface_reset.reset
			read      => mm_interconnect_0_the_altpll_pll_slave_read,      --             pll_slave.read
			write     => mm_interconnect_0_the_altpll_pll_slave_write,     --                      .write
			address   => mm_interconnect_0_the_altpll_pll_slave_address,   --                      .address
			readdata  => mm_interconnect_0_the_altpll_pll_slave_readdata,  --                      .readdata
			writedata => mm_interconnect_0_the_altpll_pll_slave_writedata, --                      .writedata
			c0        => the_altpll_c0_clk,                                --                    c0.clk
			c1        => clk_sdram_clk,                                    --                    c1.clk
			areset    => the_altpll_areset_export,                         --        areset_conduit.export
			locked    => the_altpll_locked_export,                         --        locked_conduit.export
			phasedone => the_altpll_phasedone_export                       --     phasedone_conduit.export
		);

	the_jtag_uart : component QD1_the_jtag_uart
		port map (
			clk            => clk_clk,                                                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                          --             reset.reset_n
			av_chipselect  => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_receiver_irq(0)                                   --               irq.irq
		);

	the_master : component QD1_the_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                         --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,         --    clk_reset.reset
			master_address       => the_master_master_address,       --       master.address
			master_readdata      => the_master_master_readdata,      --             .readdata
			master_read          => the_master_master_read,          --             .read
			master_write         => the_master_master_write,         --             .write
			master_writedata     => the_master_master_writedata,     --             .writedata
			master_waitrequest   => the_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => the_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => the_master_master_byteenable,    --             .byteenable
			master_reset_reset   => open                             -- master_reset.reset
		);

	the_memory_mapped_reset : component memory_mapped_reset
		generic map (
			ADDR_WIDTH    => 2,
			REGISTER_SIZE => 32
		)
		port map (
			clk               => clk_clk,                                                              --        clock.clk
			reset             => rst_controller_002_reset_out_reset,                                   --        reset.reset
			avm_address       => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_address,       -- avalon_slave.address
			avm_readdata      => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_readdata,      --             .readdata
			avm_readdatavalid => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_readdatavalid, --             .readdatavalid
			avm_read          => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_read,          --             .read
			avm_write         => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_write,         --             .write
			avm_writedata     => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_writedata,     --             .writedata
			reset_out         => the_memory_mapped_reset_reset_source_reset                            -- reset_source.reset
		);

	the_mm_clock_crossing_bridge : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 31,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk_clk,                                                         --   m0_clk.clk
			m0_reset         => rst_controller_002_reset_out_reset,                              -- m0_reset.reset
			s0_clk           => the_altpll_c0_clk,                                               --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset,                              -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_address,       --         .address
			s0_write         => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_write,         --         .write
			s0_read          => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => the_mm_clock_crossing_bridge_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => the_mm_clock_crossing_bridge_m0_readdata,                        --         .readdata
			m0_readdatavalid => the_mm_clock_crossing_bridge_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => the_mm_clock_crossing_bridge_m0_burstcount,                      --         .burstcount
			m0_writedata     => the_mm_clock_crossing_bridge_m0_writedata,                       --         .writedata
			m0_address       => the_mm_clock_crossing_bridge_m0_address,                         --         .address
			m0_write         => the_mm_clock_crossing_bridge_m0_write,                           --         .write
			m0_read          => the_mm_clock_crossing_bridge_m0_read,                            --         .read
			m0_byteenable    => the_mm_clock_crossing_bridge_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => the_mm_clock_crossing_bridge_m0_debugaccess                      --         .debugaccess
		);

	the_onchip_memory2 : component QD1_the_onchip_memory2
		port map (
			clk         => the_altpll_c0_clk,                                  --   clk1.clk
			address     => mm_interconnect_1_the_onchip_memory2_s1_address,    --     s1.address
			clken       => mm_interconnect_1_the_onchip_memory2_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_the_onchip_memory2_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_the_onchip_memory2_s1_write,      --       .write
			readdata    => mm_interconnect_1_the_onchip_memory2_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_the_onchip_memory2_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_the_onchip_memory2_s1_byteenable, --       .byteenable
			reset       => rst_controller_001_reset_out_reset,                 -- reset1.reset
			reset_req   => rst_controller_001_reset_out_reset_req,             --       .reset_req
			address2    => mm_interconnect_0_the_onchip_memory2_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_the_onchip_memory2_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_the_onchip_memory2_s2_clken,      --       .clken
			write2      => mm_interconnect_0_the_onchip_memory2_s2_write,      --       .write
			readdata2   => mm_interconnect_0_the_onchip_memory2_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_the_onchip_memory2_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_the_onchip_memory2_s2_byteenable, --       .byteenable
			clk2        => the_altpll_c0_clk,                                  --   clk2.clk
			reset2      => rst_controller_001_reset_out_reset,                 -- reset2.reset
			reset_req2  => rst_controller_001_reset_out_reset_req              --       .reset_req
		);

	the_orca_timer : component orca_timer
		generic map (
			TIMER_WIDTH => 32
		)
		port map (
			clk             => the_altpll_c0_clk,                              --           clock.clk
			reset           => rst_controller_001_reset_out_reset,             --           reset.reset
			timer_value     => the_orca_timer_timer_interface_value,           -- Timer_Interface.value
			timer_interrupt => the_orca_timer_timer_interface_interrupt,       --                .interrupt
			slave_ARADDR    => mm_interconnect_0_the_orca_timer_slave_araddr,  --           slave.araddr
			slave_ARPROT    => mm_interconnect_0_the_orca_timer_slave_arprot,  --                .arprot
			slave_ARVALID   => mm_interconnect_0_the_orca_timer_slave_arvalid, --                .arvalid
			slave_ARREADY   => mm_interconnect_0_the_orca_timer_slave_arready, --                .arready
			slave_RDATA     => mm_interconnect_0_the_orca_timer_slave_rdata,   --                .rdata
			slave_RVALID    => mm_interconnect_0_the_orca_timer_slave_rvalid,  --                .rvalid
			slave_RREADY    => mm_interconnect_0_the_orca_timer_slave_rready,  --                .rready
			slave_AWADDR    => mm_interconnect_0_the_orca_timer_slave_awaddr,  --                .awaddr
			slave_AWPROT    => mm_interconnect_0_the_orca_timer_slave_awprot,  --                .awprot
			slave_AWVALID   => mm_interconnect_0_the_orca_timer_slave_awvalid, --                .awvalid
			slave_AWREADY   => mm_interconnect_0_the_orca_timer_slave_awready, --                .awready
			slave_WDATA     => mm_interconnect_0_the_orca_timer_slave_wdata,   --                .wdata
			slave_WSTRB     => mm_interconnect_0_the_orca_timer_slave_wstrb,   --                .wstrb
			slave_WVALID    => mm_interconnect_0_the_orca_timer_slave_wvalid,  --                .wvalid
			slave_WREADY    => mm_interconnect_0_the_orca_timer_slave_wready,  --                .wready
			slave_BVALID    => mm_interconnect_0_the_orca_timer_slave_bvalid,  --                .bvalid
			slave_BREADY    => mm_interconnect_0_the_orca_timer_slave_bready,  --                .bready
			slave_BRESP     => mm_interconnect_0_the_orca_timer_slave_bresp,   --                .bresp
			slave_RRESP     => mm_interconnect_0_the_orca_timer_slave_rresp,   --                .rresp
			slave_AWLOCK    => "00",                                           --     (terminated)
			slave_ARCACHE   => "0000",                                         --     (terminated)
			slave_ARID      => "0000",                                         --     (terminated)
			slave_ARLEN     => "0000",                                         --     (terminated)
			slave_ARLOCK    => "00",                                           --     (terminated)
			slave_ARSIZE    => "000",                                          --     (terminated)
			slave_ARBURST   => "00",                                           --     (terminated)
			slave_AWBURST   => "00",                                           --     (terminated)
			slave_AWCACHE   => "0000",                                         --     (terminated)
			slave_AWID      => "0000",                                         --     (terminated)
			slave_AWLEN     => "0000",                                         --     (terminated)
			slave_AWSIZE    => "000",                                          --     (terminated)
			slave_BID       => open,                                           --     (terminated)
			slave_RID       => open,                                           --     (terminated)
			slave_RLAST     => open,                                           --     (terminated)
			slave_WID       => "0000",                                         --     (terminated)
			slave_WLAST     => '0'                                             --     (terminated)
		);

	the_vectorblox_orca : component ORCA
		generic map (
			REGISTER_SIZE                => 32,
			RESET_VECTOR                 => "00000000000000000000000000000000",
			ENABLE_EXCEPTIONS            => 1,
			INTERRUPT_VECTOR             => "00000000000000000000000000000100",
			ENABLE_EXT_INTERRUPTS        => 1,
			NUM_EXT_INTERRUPTS           => 32,
			MAX_IFETCHES_IN_FLIGHT       => 1,
			BTB_ENTRIES                  => 16,
			MULTIPLY_ENABLE              => 1,
			SHIFTER_MAX_CYCLES           => 1,
			DIVIDE_ENABLE                => 1,
			PIPELINE_STAGES              => 4,
			VCP_ENABLE                   => 0,
			POWER_OPTIMIZED              => 0,
			FAMILY                       => "ALTERA",
			INSTRUCTION_REQUEST_REGISTER => 0,
			INSTRUCTION_RETURN_REGISTER  => 0,
			DATA_REQUEST_REGISTER        => 1,
			DATA_RETURN_REGISTER         => 0,
			LOG2_BURSTLENGTH             => 4,
			AXI_ID_WIDTH                 => 2,
			AVALON_AUX                   => 1,
			LMB_AUX                      => 0,
			WISHBONE_AUX                 => 0,
			ICACHE_SIZE                  => 0,
			ICACHE_LINE_SIZE             => 32,
			ICACHE_EXTERNAL_WIDTH        => 32,
			IC_REQUEST_REGISTER          => 1,
			IC_RETURN_REGISTER           => 0,
			DCACHE_SIZE                  => 0,
			DCACHE_WRITEBACK             => 1,
			DCACHE_LINE_SIZE             => 32,
			DCACHE_EXTERNAL_WIDTH        => 32,
			DC_REQUEST_REGISTER          => 1,
			DC_RETURN_REGISTER           => 0,
			UC_MEMORY_REGIONS            => 0,
			UMR0_ADDR_BASE               => "00000000000000000000000000000000",
			UMR0_ADDR_LAST               => "00000000000000000000000000000000",
			IUC_REQUEST_REGISTER         => 1,
			IUC_RETURN_REGISTER          => 0,
			DUC_REQUEST_REGISTER         => 2,
			DUC_RETURN_REGISTER          => 1,
			AUX_MEMORY_REGIONS           => 1,
			AMR0_ADDR_BASE               => "00000000000000000000000000000000",
			AMR0_ADDR_LAST               => "11111111111111111111111111111111",
			IAUX_REQUEST_REGISTER        => 0,
			IAUX_RETURN_REGISTER         => 0,
			DAUX_REQUEST_REGISTER        => 0,
			DAUX_RETURN_REGISTER         => 0
		)
		port map (
			clk                           => the_altpll_c0_clk,                             --             clock.clk
			reset                         => rst_controller_003_reset_out_reset,            --             reset.reset
			avm_data_address              => the_vectorblox_orca_data_address,              --              data.address
			avm_data_byteenable           => the_vectorblox_orca_data_byteenable,           --                  .byteenable
			avm_data_read                 => the_vectorblox_orca_data_read,                 --                  .read
			avm_data_readdata             => the_vectorblox_orca_data_readdata,             --                  .readdata
			avm_data_write                => the_vectorblox_orca_data_write,                --                  .write
			avm_data_writedata            => the_vectorblox_orca_data_writedata,            --                  .writedata
			avm_data_waitrequest          => the_vectorblox_orca_data_waitrequest,          --                  .waitrequest
			avm_data_readdatavalid        => the_vectorblox_orca_data_readdatavalid,        --                  .readdatavalid
			avm_instruction_address       => the_vectorblox_orca_instruction_address,       --       instruction.address
			avm_instruction_read          => the_vectorblox_orca_instruction_read,          --                  .read
			avm_instruction_readdata      => the_vectorblox_orca_instruction_readdata,      --                  .readdata
			avm_instruction_waitrequest   => the_vectorblox_orca_instruction_waitrequest,   --                  .waitrequest
			avm_instruction_readdatavalid => the_vectorblox_orca_instruction_readdatavalid, --                  .readdatavalid
			timer_value                   => the_orca_timer_timer_interface_value,          --   Timer_Interface.value
			timer_interrupt               => the_orca_timer_timer_interface_interrupt,      --                  .interrupt
			global_interrupts             => the_vectorblox_orca_global_interrupts_irq,     -- global_interrupts.irq
			DUC_ARADDR                    => open,                                          --       (terminated)
			DUC_ARBURST                   => open,                                          --       (terminated)
			DUC_ARCACHE                   => open,                                          --       (terminated)
			DUC_ARID                      => open,                                          --       (terminated)
			DUC_ARLEN                     => open,                                          --       (terminated)
			DUC_ARLOCK                    => open,                                          --       (terminated)
			DUC_ARPROT                    => open,                                          --       (terminated)
			DUC_ARREADY                   => '0',                                           --       (terminated)
			DUC_ARSIZE                    => open,                                          --       (terminated)
			DUC_ARVALID                   => open,                                          --       (terminated)
			DUC_AWADDR                    => open,                                          --       (terminated)
			DUC_AWBURST                   => open,                                          --       (terminated)
			DUC_AWCACHE                   => open,                                          --       (terminated)
			DUC_AWID                      => open,                                          --       (terminated)
			DUC_AWLEN                     => open,                                          --       (terminated)
			DUC_AWLOCK                    => open,                                          --       (terminated)
			DUC_AWPROT                    => open,                                          --       (terminated)
			DUC_AWREADY                   => '0',                                           --       (terminated)
			DUC_AWSIZE                    => open,                                          --       (terminated)
			DUC_AWVALID                   => open,                                          --       (terminated)
			DUC_BID                       => "00",                                          --       (terminated)
			DUC_BREADY                    => open,                                          --       (terminated)
			DUC_BRESP                     => "00",                                          --       (terminated)
			DUC_BVALID                    => '0',                                           --       (terminated)
			DUC_RDATA                     => "00000000000000000000000000000000",            --       (terminated)
			DUC_RID                       => "00",                                          --       (terminated)
			DUC_RLAST                     => '0',                                           --       (terminated)
			DUC_RREADY                    => open,                                          --       (terminated)
			DUC_RRESP                     => "00",                                          --       (terminated)
			DUC_RVALID                    => '0',                                           --       (terminated)
			DUC_WDATA                     => open,                                          --       (terminated)
			DUC_WID                       => open,                                          --       (terminated)
			DUC_WLAST                     => open,                                          --       (terminated)
			DUC_WREADY                    => '0',                                           --       (terminated)
			DUC_WSTRB                     => open,                                          --       (terminated)
			DUC_WVALID                    => open,                                          --       (terminated)
			IUC_ARADDR                    => open,                                          --       (terminated)
			IUC_ARBURST                   => open,                                          --       (terminated)
			IUC_ARCACHE                   => open,                                          --       (terminated)
			IUC_ARID                      => open,                                          --       (terminated)
			IUC_ARLEN                     => open,                                          --       (terminated)
			IUC_ARLOCK                    => open,                                          --       (terminated)
			IUC_ARPROT                    => open,                                          --       (terminated)
			IUC_ARREADY                   => '0',                                           --       (terminated)
			IUC_ARSIZE                    => open,                                          --       (terminated)
			IUC_ARVALID                   => open,                                          --       (terminated)
			IUC_AWADDR                    => open,                                          --       (terminated)
			IUC_AWBURST                   => open,                                          --       (terminated)
			IUC_AWCACHE                   => open,                                          --       (terminated)
			IUC_AWID                      => open,                                          --       (terminated)
			IUC_AWLEN                     => open,                                          --       (terminated)
			IUC_AWLOCK                    => open,                                          --       (terminated)
			IUC_AWPROT                    => open,                                          --       (terminated)
			IUC_AWREADY                   => '0',                                           --       (terminated)
			IUC_AWSIZE                    => open,                                          --       (terminated)
			IUC_AWVALID                   => open,                                          --       (terminated)
			IUC_BID                       => "00",                                          --       (terminated)
			IUC_BREADY                    => open,                                          --       (terminated)
			IUC_BRESP                     => "00",                                          --       (terminated)
			IUC_BVALID                    => '0',                                           --       (terminated)
			IUC_RDATA                     => "00000000000000000000000000000000",            --       (terminated)
			IUC_RID                       => "00",                                          --       (terminated)
			IUC_RLAST                     => '0',                                           --       (terminated)
			IUC_RREADY                    => open,                                          --       (terminated)
			IUC_RRESP                     => "00",                                          --       (terminated)
			IUC_RVALID                    => '0',                                           --       (terminated)
			IUC_WDATA                     => open,                                          --       (terminated)
			IUC_WID                       => open,                                          --       (terminated)
			IUC_WLAST                     => open,                                          --       (terminated)
			IUC_WREADY                    => '0',                                           --       (terminated)
			IUC_WSTRB                     => open,                                          --       (terminated)
			IUC_WVALID                    => open,                                          --       (terminated)
			IC_ARADDR                     => open,                                          --       (terminated)
			IC_ARBURST                    => open,                                          --       (terminated)
			IC_ARCACHE                    => open,                                          --       (terminated)
			IC_ARID                       => open,                                          --       (terminated)
			IC_ARLEN                      => open,                                          --       (terminated)
			IC_ARLOCK                     => open,                                          --       (terminated)
			IC_ARPROT                     => open,                                          --       (terminated)
			IC_ARREADY                    => '0',                                           --       (terminated)
			IC_ARSIZE                     => open,                                          --       (terminated)
			IC_ARVALID                    => open,                                          --       (terminated)
			IC_AWADDR                     => open,                                          --       (terminated)
			IC_AWBURST                    => open,                                          --       (terminated)
			IC_AWCACHE                    => open,                                          --       (terminated)
			IC_AWID                       => open,                                          --       (terminated)
			IC_AWLEN                      => open,                                          --       (terminated)
			IC_AWLOCK                     => open,                                          --       (terminated)
			IC_AWPROT                     => open,                                          --       (terminated)
			IC_AWREADY                    => '0',                                           --       (terminated)
			IC_AWSIZE                     => open,                                          --       (terminated)
			IC_AWVALID                    => open,                                          --       (terminated)
			IC_BID                        => "00",                                          --       (terminated)
			IC_BREADY                     => open,                                          --       (terminated)
			IC_BRESP                      => "00",                                          --       (terminated)
			IC_BVALID                     => '0',                                           --       (terminated)
			IC_RDATA                      => "00000000000000000000000000000000",            --       (terminated)
			IC_RID                        => "00",                                          --       (terminated)
			IC_RLAST                      => '0',                                           --       (terminated)
			IC_RREADY                     => open,                                          --       (terminated)
			IC_RRESP                      => "00",                                          --       (terminated)
			IC_RVALID                     => '0',                                           --       (terminated)
			IC_WDATA                      => open,                                          --       (terminated)
			IC_WID                        => open,                                          --       (terminated)
			IC_WLAST                      => open,                                          --       (terminated)
			IC_WREADY                     => '0',                                           --       (terminated)
			IC_WSTRB                      => open,                                          --       (terminated)
			IC_WVALID                     => open,                                          --       (terminated)
			DC_ARADDR                     => open,                                          --       (terminated)
			DC_ARBURST                    => open,                                          --       (terminated)
			DC_ARCACHE                    => open,                                          --       (terminated)
			DC_ARID                       => open,                                          --       (terminated)
			DC_ARLEN                      => open,                                          --       (terminated)
			DC_ARLOCK                     => open,                                          --       (terminated)
			DC_ARPROT                     => open,                                          --       (terminated)
			DC_ARREADY                    => '0',                                           --       (terminated)
			DC_ARSIZE                     => open,                                          --       (terminated)
			DC_ARVALID                    => open,                                          --       (terminated)
			DC_AWADDR                     => open,                                          --       (terminated)
			DC_AWBURST                    => open,                                          --       (terminated)
			DC_AWCACHE                    => open,                                          --       (terminated)
			DC_AWID                       => open,                                          --       (terminated)
			DC_AWLEN                      => open,                                          --       (terminated)
			DC_AWLOCK                     => open,                                          --       (terminated)
			DC_AWPROT                     => open,                                          --       (terminated)
			DC_AWREADY                    => '0',                                           --       (terminated)
			DC_AWSIZE                     => open,                                          --       (terminated)
			DC_AWVALID                    => open,                                          --       (terminated)
			DC_BID                        => "00",                                          --       (terminated)
			DC_BREADY                     => open,                                          --       (terminated)
			DC_BRESP                      => "00",                                          --       (terminated)
			DC_BVALID                     => '0',                                           --       (terminated)
			DC_RDATA                      => "00000000000000000000000000000000",            --       (terminated)
			DC_RID                        => "00",                                          --       (terminated)
			DC_RLAST                      => '0',                                           --       (terminated)
			DC_RREADY                     => open,                                          --       (terminated)
			DC_RRESP                      => "00",                                          --       (terminated)
			DC_RVALID                     => '0',                                           --       (terminated)
			DC_WDATA                      => open,                                          --       (terminated)
			DC_WID                        => open,                                          --       (terminated)
			DC_WLAST                      => open,                                          --       (terminated)
			DC_WREADY                     => '0',                                           --       (terminated)
			DC_WSTRB                      => open,                                          --       (terminated)
			DC_WVALID                     => open,                                          --       (terminated)
			vcp_data0                     => open,                                          --       (terminated)
			vcp_data1                     => open,                                          --       (terminated)
			vcp_data2                     => open,                                          --       (terminated)
			vcp_instruction               => open,                                          --       (terminated)
			vcp_valid_instr               => open,                                          --       (terminated)
			vcp_ready                     => '0',                                           --       (terminated)
			vcp_illegal                   => '0',                                           --       (terminated)
			vcp_writeback_data            => "00000000000000000000000000000000",            --       (terminated)
			vcp_writeback_en              => '0',                                           --       (terminated)
			vcp_alu_data1                 => "00000000000000000000000000000000",            --       (terminated)
			vcp_alu_data2                 => "00000000000000000000000000000000",            --       (terminated)
			vcp_alu_source_valid          => '0',                                           --       (terminated)
			vcp_alu_result                => open,                                          --       (terminated)
			vcp_alu_result_valid          => open,                                          --       (terminated)
			data_ADR_O                    => open,                                          --       (terminated)
			data_DAT_I                    => "00000000000000000000000000000000",            --       (terminated)
			data_DAT_O                    => open,                                          --       (terminated)
			data_WE_O                     => open,                                          --       (terminated)
			data_SEL_O                    => open,                                          --       (terminated)
			data_STB_O                    => open,                                          --       (terminated)
			data_ACK_I                    => '0',                                           --       (terminated)
			data_CYC_O                    => open,                                          --       (terminated)
			data_CTI_O                    => open,                                          --       (terminated)
			data_STALL_I                  => '0',                                           --       (terminated)
			instr_ADR_O                   => open,                                          --       (terminated)
			instr_DAT_I                   => "00000000000000000000000000000000",            --       (terminated)
			instr_STB_O                   => open,                                          --       (terminated)
			instr_ACK_I                   => '0',                                           --       (terminated)
			instr_CYC_O                   => open,                                          --       (terminated)
			instr_CTI_O                   => open,                                          --       (terminated)
			instr_STALL_I                 => '0',                                           --       (terminated)
			ILMB_Addr                     => open,                                          --       (terminated)
			ILMB_Byte_Enable              => open,                                          --       (terminated)
			ILMB_Data_Write               => open,                                          --       (terminated)
			ILMB_AS                       => open,                                          --       (terminated)
			ILMB_Read_Strobe              => open,                                          --       (terminated)
			ILMB_Write_Strobe             => open,                                          --       (terminated)
			ILMB_Data_Read                => "00000000000000000000000000000000",            --       (terminated)
			ILMB_Ready                    => '0',                                           --       (terminated)
			ILMB_Wait                     => '0',                                           --       (terminated)
			ILMB_CE                       => '0',                                           --       (terminated)
			ILMB_UE                       => '0',                                           --       (terminated)
			DLMB_Addr                     => open,                                          --       (terminated)
			DLMB_Byte_Enable              => open,                                          --       (terminated)
			DLMB_Data_Write               => open,                                          --       (terminated)
			DLMB_AS                       => open,                                          --       (terminated)
			DLMB_Read_Strobe              => open,                                          --       (terminated)
			DLMB_Write_Strobe             => open,                                          --       (terminated)
			DLMB_Data_Read                => "00000000000000000000000000000000",            --       (terminated)
			DLMB_Ready                    => '0',                                           --       (terminated)
			DLMB_Wait                     => '0',                                           --       (terminated)
			DLMB_CE                       => '0',                                           --       (terminated)
			DLMB_UE                       => '0'                                            --       (terminated)
		);

	mm_interconnect_0 : component QD1_mm_interconnect_0
		port map (
			the_orca_timer_slave_awaddr                                       => mm_interconnect_0_the_orca_timer_slave_awaddr,                        --                                        the_orca_timer_slave.awaddr
			the_orca_timer_slave_awprot                                       => mm_interconnect_0_the_orca_timer_slave_awprot,                        --                                                            .awprot
			the_orca_timer_slave_awvalid                                      => mm_interconnect_0_the_orca_timer_slave_awvalid,                       --                                                            .awvalid
			the_orca_timer_slave_awready                                      => mm_interconnect_0_the_orca_timer_slave_awready,                       --                                                            .awready
			the_orca_timer_slave_wdata                                        => mm_interconnect_0_the_orca_timer_slave_wdata,                         --                                                            .wdata
			the_orca_timer_slave_wstrb                                        => mm_interconnect_0_the_orca_timer_slave_wstrb,                         --                                                            .wstrb
			the_orca_timer_slave_wvalid                                       => mm_interconnect_0_the_orca_timer_slave_wvalid,                        --                                                            .wvalid
			the_orca_timer_slave_wready                                       => mm_interconnect_0_the_orca_timer_slave_wready,                        --                                                            .wready
			the_orca_timer_slave_bresp                                        => mm_interconnect_0_the_orca_timer_slave_bresp,                         --                                                            .bresp
			the_orca_timer_slave_bvalid                                       => mm_interconnect_0_the_orca_timer_slave_bvalid,                        --                                                            .bvalid
			the_orca_timer_slave_bready                                       => mm_interconnect_0_the_orca_timer_slave_bready,                        --                                                            .bready
			the_orca_timer_slave_araddr                                       => mm_interconnect_0_the_orca_timer_slave_araddr,                        --                                                            .araddr
			the_orca_timer_slave_arprot                                       => mm_interconnect_0_the_orca_timer_slave_arprot,                        --                                                            .arprot
			the_orca_timer_slave_arvalid                                      => mm_interconnect_0_the_orca_timer_slave_arvalid,                       --                                                            .arvalid
			the_orca_timer_slave_arready                                      => mm_interconnect_0_the_orca_timer_slave_arready,                       --                                                            .arready
			the_orca_timer_slave_rdata                                        => mm_interconnect_0_the_orca_timer_slave_rdata,                         --                                                            .rdata
			the_orca_timer_slave_rresp                                        => mm_interconnect_0_the_orca_timer_slave_rresp,                         --                                                            .rresp
			the_orca_timer_slave_rvalid                                       => mm_interconnect_0_the_orca_timer_slave_rvalid,                        --                                                            .rvalid
			the_orca_timer_slave_rready                                       => mm_interconnect_0_the_orca_timer_slave_rready,                        --                                                            .rready
			the_altpll_c0_clk                                                 => the_altpll_c0_clk,                                                    --                                               the_altpll_c0.clk
			the_clk_clk_clk                                                   => clk_clk,                                                              --                                                 the_clk_clk.clk
			the_altpll_inclk_interface_reset_reset_bridge_in_reset_reset      => rst_controller_002_reset_out_reset,                                   --      the_altpll_inclk_interface_reset_reset_bridge_in_reset.reset
			the_jtag_uart_reset_reset_bridge_in_reset_reset                   => rst_controller_reset_out_reset,                                       --                   the_jtag_uart_reset_reset_bridge_in_reset.reset
			the_master_clk_reset_reset_bridge_in_reset_reset                  => rst_controller_002_reset_out_reset,                                   --                  the_master_clk_reset_reset_bridge_in_reset.reset
			the_mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                   -- the_mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset.reset
			the_vectorblox_orca_reset_reset_bridge_in_reset_reset             => rst_controller_003_reset_out_reset,                                   --             the_vectorblox_orca_reset_reset_bridge_in_reset.reset
			the_master_master_address                                         => the_master_master_address,                                            --                                           the_master_master.address
			the_master_master_waitrequest                                     => the_master_master_waitrequest,                                        --                                                            .waitrequest
			the_master_master_byteenable                                      => the_master_master_byteenable,                                         --                                                            .byteenable
			the_master_master_read                                            => the_master_master_read,                                               --                                                            .read
			the_master_master_readdata                                        => the_master_master_readdata,                                           --                                                            .readdata
			the_master_master_readdatavalid                                   => the_master_master_readdatavalid,                                      --                                                            .readdatavalid
			the_master_master_write                                           => the_master_master_write,                                              --                                                            .write
			the_master_master_writedata                                       => the_master_master_writedata,                                          --                                                            .writedata
			the_mm_clock_crossing_bridge_m0_address                           => the_mm_clock_crossing_bridge_m0_address,                              --                             the_mm_clock_crossing_bridge_m0.address
			the_mm_clock_crossing_bridge_m0_waitrequest                       => the_mm_clock_crossing_bridge_m0_waitrequest,                          --                                                            .waitrequest
			the_mm_clock_crossing_bridge_m0_burstcount                        => the_mm_clock_crossing_bridge_m0_burstcount,                           --                                                            .burstcount
			the_mm_clock_crossing_bridge_m0_byteenable                        => the_mm_clock_crossing_bridge_m0_byteenable,                           --                                                            .byteenable
			the_mm_clock_crossing_bridge_m0_read                              => the_mm_clock_crossing_bridge_m0_read,                                 --                                                            .read
			the_mm_clock_crossing_bridge_m0_readdata                          => the_mm_clock_crossing_bridge_m0_readdata,                             --                                                            .readdata
			the_mm_clock_crossing_bridge_m0_readdatavalid                     => the_mm_clock_crossing_bridge_m0_readdatavalid,                        --                                                            .readdatavalid
			the_mm_clock_crossing_bridge_m0_write                             => the_mm_clock_crossing_bridge_m0_write,                                --                                                            .write
			the_mm_clock_crossing_bridge_m0_writedata                         => the_mm_clock_crossing_bridge_m0_writedata,                            --                                                            .writedata
			the_mm_clock_crossing_bridge_m0_debugaccess                       => the_mm_clock_crossing_bridge_m0_debugaccess,                          --                                                            .debugaccess
			the_vectorblox_orca_data_address                                  => the_vectorblox_orca_data_address,                                     --                                    the_vectorblox_orca_data.address
			the_vectorblox_orca_data_waitrequest                              => the_vectorblox_orca_data_waitrequest,                                 --                                                            .waitrequest
			the_vectorblox_orca_data_byteenable                               => the_vectorblox_orca_data_byteenable,                                  --                                                            .byteenable
			the_vectorblox_orca_data_read                                     => the_vectorblox_orca_data_read,                                        --                                                            .read
			the_vectorblox_orca_data_readdata                                 => the_vectorblox_orca_data_readdata,                                    --                                                            .readdata
			the_vectorblox_orca_data_readdatavalid                            => the_vectorblox_orca_data_readdatavalid,                               --                                                            .readdatavalid
			the_vectorblox_orca_data_write                                    => the_vectorblox_orca_data_write,                                       --                                                            .write
			the_vectorblox_orca_data_writedata                                => the_vectorblox_orca_data_writedata,                                   --                                                            .writedata
			button_pio_s1_address                                             => mm_interconnect_0_button_pio_s1_address,                              --                                               button_pio_s1.address
			button_pio_s1_write                                               => mm_interconnect_0_button_pio_s1_write,                                --                                                            .write
			button_pio_s1_readdata                                            => mm_interconnect_0_button_pio_s1_readdata,                             --                                                            .readdata
			button_pio_s1_writedata                                           => mm_interconnect_0_button_pio_s1_writedata,                            --                                                            .writedata
			button_pio_s1_chipselect                                          => mm_interconnect_0_button_pio_s1_chipselect,                           --                                                            .chipselect
			led_pio_s1_address                                                => mm_interconnect_0_led_pio_s1_address,                                 --                                                  led_pio_s1.address
			led_pio_s1_write                                                  => mm_interconnect_0_led_pio_s1_write,                                   --                                                            .write
			led_pio_s1_readdata                                               => mm_interconnect_0_led_pio_s1_readdata,                                --                                                            .readdata
			led_pio_s1_writedata                                              => mm_interconnect_0_led_pio_s1_writedata,                               --                                                            .writedata
			led_pio_s1_chipselect                                             => mm_interconnect_0_led_pio_s1_chipselect,                              --                                                            .chipselect
			sdram_s1_address                                                  => mm_interconnect_0_sdram_s1_address,                                   --                                                    sdram_s1.address
			sdram_s1_write                                                    => mm_interconnect_0_sdram_s1_write,                                     --                                                            .write
			sdram_s1_read                                                     => mm_interconnect_0_sdram_s1_read,                                      --                                                            .read
			sdram_s1_readdata                                                 => mm_interconnect_0_sdram_s1_readdata,                                  --                                                            .readdata
			sdram_s1_writedata                                                => mm_interconnect_0_sdram_s1_writedata,                                 --                                                            .writedata
			sdram_s1_byteenable                                               => mm_interconnect_0_sdram_s1_byteenable,                                --                                                            .byteenable
			sdram_s1_readdatavalid                                            => mm_interconnect_0_sdram_s1_readdatavalid,                             --                                                            .readdatavalid
			sdram_s1_waitrequest                                              => mm_interconnect_0_sdram_s1_waitrequest,                               --                                                            .waitrequest
			sdram_s1_chipselect                                               => mm_interconnect_0_sdram_s1_chipselect,                                --                                                            .chipselect
			switch_pio_s1_address                                             => mm_interconnect_0_switch_pio_s1_address,                              --                                               switch_pio_s1.address
			switch_pio_s1_readdata                                            => mm_interconnect_0_switch_pio_s1_readdata,                             --                                                            .readdata
			the_altpll_pll_slave_address                                      => mm_interconnect_0_the_altpll_pll_slave_address,                       --                                        the_altpll_pll_slave.address
			the_altpll_pll_slave_write                                        => mm_interconnect_0_the_altpll_pll_slave_write,                         --                                                            .write
			the_altpll_pll_slave_read                                         => mm_interconnect_0_the_altpll_pll_slave_read,                          --                                                            .read
			the_altpll_pll_slave_readdata                                     => mm_interconnect_0_the_altpll_pll_slave_readdata,                      --                                                            .readdata
			the_altpll_pll_slave_writedata                                    => mm_interconnect_0_the_altpll_pll_slave_writedata,                     --                                                            .writedata
			the_jtag_uart_avalon_jtag_slave_address                           => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_address,            --                             the_jtag_uart_avalon_jtag_slave.address
			the_jtag_uart_avalon_jtag_slave_write                             => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write,              --                                                            .write
			the_jtag_uart_avalon_jtag_slave_read                              => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read,               --                                                            .read
			the_jtag_uart_avalon_jtag_slave_readdata                          => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_readdata,           --                                                            .readdata
			the_jtag_uart_avalon_jtag_slave_writedata                         => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_writedata,          --                                                            .writedata
			the_jtag_uart_avalon_jtag_slave_waitrequest                       => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_waitrequest,        --                                                            .waitrequest
			the_jtag_uart_avalon_jtag_slave_chipselect                        => mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_chipselect,         --                                                            .chipselect
			the_memory_mapped_reset_avalon_slave_address                      => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_address,       --                        the_memory_mapped_reset_avalon_slave.address
			the_memory_mapped_reset_avalon_slave_write                        => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_write,         --                                                            .write
			the_memory_mapped_reset_avalon_slave_read                         => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_read,          --                                                            .read
			the_memory_mapped_reset_avalon_slave_readdata                     => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_readdata,      --                                                            .readdata
			the_memory_mapped_reset_avalon_slave_writedata                    => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_writedata,     --                                                            .writedata
			the_memory_mapped_reset_avalon_slave_readdatavalid                => mm_interconnect_0_the_memory_mapped_reset_avalon_slave_readdatavalid, --                                                            .readdatavalid
			the_mm_clock_crossing_bridge_s0_address                           => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_address,            --                             the_mm_clock_crossing_bridge_s0.address
			the_mm_clock_crossing_bridge_s0_write                             => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_write,              --                                                            .write
			the_mm_clock_crossing_bridge_s0_read                              => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_read,               --                                                            .read
			the_mm_clock_crossing_bridge_s0_readdata                          => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_readdata,           --                                                            .readdata
			the_mm_clock_crossing_bridge_s0_writedata                         => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_writedata,          --                                                            .writedata
			the_mm_clock_crossing_bridge_s0_burstcount                        => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_burstcount,         --                                                            .burstcount
			the_mm_clock_crossing_bridge_s0_byteenable                        => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_byteenable,         --                                                            .byteenable
			the_mm_clock_crossing_bridge_s0_readdatavalid                     => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_readdatavalid,      --                                                            .readdatavalid
			the_mm_clock_crossing_bridge_s0_waitrequest                       => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_waitrequest,        --                                                            .waitrequest
			the_mm_clock_crossing_bridge_s0_debugaccess                       => mm_interconnect_0_the_mm_clock_crossing_bridge_s0_debugaccess,        --                                                            .debugaccess
			the_onchip_memory2_s2_address                                     => mm_interconnect_0_the_onchip_memory2_s2_address,                      --                                       the_onchip_memory2_s2.address
			the_onchip_memory2_s2_write                                       => mm_interconnect_0_the_onchip_memory2_s2_write,                        --                                                            .write
			the_onchip_memory2_s2_readdata                                    => mm_interconnect_0_the_onchip_memory2_s2_readdata,                     --                                                            .readdata
			the_onchip_memory2_s2_writedata                                   => mm_interconnect_0_the_onchip_memory2_s2_writedata,                    --                                                            .writedata
			the_onchip_memory2_s2_byteenable                                  => mm_interconnect_0_the_onchip_memory2_s2_byteenable,                   --                                                            .byteenable
			the_onchip_memory2_s2_chipselect                                  => mm_interconnect_0_the_onchip_memory2_s2_chipselect,                   --                                                            .chipselect
			the_onchip_memory2_s2_clken                                       => mm_interconnect_0_the_onchip_memory2_s2_clken                         --                                                            .clken
		);

	mm_interconnect_1 : component QD1_mm_interconnect_1
		port map (
			the_altpll_c0_clk                                     => the_altpll_c0_clk,                                  --                                   the_altpll_c0.clk
			the_onchip_memory2_reset1_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                 -- the_onchip_memory2_reset1_reset_bridge_in_reset.reset
			the_vectorblox_orca_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                 -- the_vectorblox_orca_reset_reset_bridge_in_reset.reset
			the_vectorblox_orca_instruction_address               => the_vectorblox_orca_instruction_address,            --                 the_vectorblox_orca_instruction.address
			the_vectorblox_orca_instruction_waitrequest           => the_vectorblox_orca_instruction_waitrequest,        --                                                .waitrequest
			the_vectorblox_orca_instruction_read                  => the_vectorblox_orca_instruction_read,               --                                                .read
			the_vectorblox_orca_instruction_readdata              => the_vectorblox_orca_instruction_readdata,           --                                                .readdata
			the_vectorblox_orca_instruction_readdatavalid         => the_vectorblox_orca_instruction_readdatavalid,      --                                                .readdatavalid
			the_onchip_memory2_s1_address                         => mm_interconnect_1_the_onchip_memory2_s1_address,    --                           the_onchip_memory2_s1.address
			the_onchip_memory2_s1_write                           => mm_interconnect_1_the_onchip_memory2_s1_write,      --                                                .write
			the_onchip_memory2_s1_readdata                        => mm_interconnect_1_the_onchip_memory2_s1_readdata,   --                                                .readdata
			the_onchip_memory2_s1_writedata                       => mm_interconnect_1_the_onchip_memory2_s1_writedata,  --                                                .writedata
			the_onchip_memory2_s1_byteenable                      => mm_interconnect_1_the_onchip_memory2_s1_byteenable, --                                                .byteenable
			the_onchip_memory2_s1_chipselect                      => mm_interconnect_1_the_onchip_memory2_s1_chipselect, --                                                .chipselect
			the_onchip_memory2_s1_clken                           => mm_interconnect_1_the_onchip_memory2_s1_clken       --                                                .clken
		);

	irq_mapper : component QD1_irq_mapper
		port map (
			clk           => the_altpll_c0_clk,                         --       clk.clk
			reset         => rst_controller_003_reset_out_reset,        -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,                  -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,                  -- receiver1.irq
			sender_irq    => the_vectorblox_orca_global_interrupts_irq  --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => the_altpll_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_003_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk_clk,                            --       receiver_clk.clk
			sender_clk     => the_altpll_c0_clk,                  --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_003_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	rst_controller : component qd1_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => the_memory_mapped_reset_reset_source_reset, -- reset_in1.reset
			clk            => clk_clk,                                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_001 : component qd1_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => the_altpll_c0_clk,                      --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component qd1_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component qd1_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                    -- reset_in0.reset
			reset_in1      => the_memory_mapped_reset_reset_source_reset, -- reset_in1.reset
			clk            => the_altpll_c0_clk,                          --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_the_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_button_pio_s1_write_ports_inv <= not mm_interconnect_0_button_pio_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of QD1
